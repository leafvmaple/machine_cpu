// 16 bit Adder

`ifndef _MACHINE_V_
`define _MACHINE_V_ 

`include "cpu_top.v"

module Board;

CPU cpu();

endmodule

`endif